// EECE3324 Computer Architecture
// Hw 6
// Tim Liming

// The small ALU control unit that takes the ALUop and 6-bit function code in and 
// generates 4-bit ALU_operation signal for the ALU.  

`timescale 1ns / 1ns

module ALU_control_unit(ALUop, addi, func, ALUoperation);
  
  input [1:0] ALUop;
  input addi;
  input [5:0] func;
  output reg [3:0] ALUoperation;
  
  always @ (ALUop or func) begin
    
    ALUoperation <= 4'b0000;
    
    case (ALUop)
      
      // lw & sw
      2'b00: begin ALUoperation <= 4'b0000; end
      
      // beq
      2'b01: begin ALUoperation <= 4'b0110; end
      
      // 
      2'b10: begin
        case (addi)
          1'b1: begin ALUoperation <= 4'b0000; end
          1'b0: begin
            case (func[3:0])
              // add
              4'b0000: begin ALUoperation <= 4'b0000; end
              // sub
              4'b0010: begin ALUoperation <= 4'b0110; end
              // and
              4'b0100: begin ALUoperation <= 4'b0000; end
              // or
              4'b0101: begin ALUoperation <= 4'b0001; end
              // slt
              4'b1010: begin ALUoperation <= 4'b0111; end
              default: begin ALUoperation <= 4'b0000; end
            endcase
          end
        endcase
      end
      
      // 
      2'b11: begin
        case (func[3:0])
          // sub
          4'b0010: begin ALUoperation <= 4'b0110; end
          // slt
          4'b1010: begin ALUoperation <= 4'b0111; end
          default: begin ALUoperation <= 4'b0000; end
        endcase
      end
      default: begin ALUoperation <= 4'b0000; end
    endcase
  end
  
endmodule
            
      